`timescale 1ns / 1ps

module sra8(
    input [7:0] a,    
    input [7:0] b,  
    output [7:0] out   
);

endmodule
