`timescale 1ns / 1ps

module ham32 (
    input [31:0]a,
    output [31:0]out
    );
    assign out = 0;

endmodule
