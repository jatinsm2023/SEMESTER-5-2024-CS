`timescale 1ns / 1ps

module ham8(
 
    );
endmodule
