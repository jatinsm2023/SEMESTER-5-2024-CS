`timescale 1ns / 1ps

module sl8(
    input [7:0] a,    
    input [7:0] b,  
    output [7:0] out   
);
 
endmodule
